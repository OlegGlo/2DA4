
module displaydriver();

	// === Input / Output ===	 
	
	// === Net / Reg ===
	
	// === Logic ===


endmodule
