
module adder();

	// === Input / Output ===
	
	// === Net / Reg ===
	
	// === Logic ===

endmodule
