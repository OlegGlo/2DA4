
module simpleadder(SW, HEX5);

	// === Input / Output ===
	
	// === Net / Reg ===
	
	// === Logic ===
	

endmodule
